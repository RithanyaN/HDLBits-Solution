module top_module( output one );

    assign one = 1'b1;//assign will continuously allow to update the input to the output.

endmodule
