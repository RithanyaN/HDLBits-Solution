module top_module ( 
    input p1a, p1b, p1c, p1d, p1e, p1f,
    output p1y,
    input p2a, p2b, p2c, p2d,
    output p2y );
    wire w[3:0];
    and g1(w[0],p2a,p2b);
    and g2(w[1],p2c,p2d);
    or g3(p2y,w[0],w[1]);
    and g4(w[2],p1a,p1b,p1c);
    and g5(w[3],p1d,p1e,p1f);
    or g6(p1y,w[2],w[3]);
endmodule
