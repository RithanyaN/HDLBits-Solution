module top_module( 
    input a, 
    input b, 
    output out );
    and g(out,a,b);
    //assign out = a & b;
    //assign out = a && b;
    

endmodule
