module top_module( input in, output out );
    not g(out,in);

endmodule
